// Design a 32:5 encoder using behavioral level of abstraction.

// Total output is 5 bit, input is 32 bit, and 1 bit enable

module encoder_32to5(output [4:0] out, 
                     input [31:0] in);

// truth table
/*
in[32:0] : out[4:0]
1000_0000_0000_0000_0000_0000_0000_0000 : 11111
0100_0000_0000_0000_0000_0000_0000_0000 : 11110
0010_0000_0000_0000_0000_0000_0000_0000 : 11101
0001_0000_0000_0000_0000_0000_0000_0000 : 11100
0000_1000_0000_0000_0000_0000_0000_0000 : 11011
0000_0100_0000_0000_0000_0000_0000_0000 : 11010
0000_0010_0000_0000_0000_0000_0000_0000 : 11001
0000_0001_0000_0000_0000_0000_0000_0000 : 11000
0000_0000_1000_0000_0000_0000_0000_0000 : 10111
0000_0000_0100_0000_0000_0000_0000_0000 : 10110
0000_0000_0010_0000_0000_0000_0000_0000 : 10101
0000_0000_0001_0000_0000_0000_0000_0000 : 10100
0000_0000_0000_1000_0000_0000_0000_0000 : 10011
0000_0000_0000_0100_0000_0000_0000_0000 : 10010
0000_0000_0000_0010_0000_0000_0000_0000 : 10001
0000_0000_0000_0001_0000_0000_0000_0000 : 10000
0000_0000_0000_0000_1000_0000_0000_0000 : 01111
0000_0000_0000_0000_0100_0000_0000_0000 : 01110
0000_0000_0000_0000_0010_0000_0000_0000 : 01101
0000_0000_0000_0000_0001_0000_0000_0000 : 01100
0000_0000_0000_0000_0000_1000_0000_0000 : 01011
0000_0000_0000_0000_0000_0100_0000_0000 : 01010
0000_0000_0000_0000_0000_0010_0000_0000 : 01001
0000_0000_0000_0000_0000_0001_0000_0000 : 01000
0000_0000_0000_0000_0000_0000_1000_0000 : 00111
0000_0000_0000_0000_0000_0000_0100_0000 : 00110
0000_0000_0000_0000_0000_0000_0010_0000 : 00101
0000_0000_0000_0000_0000_0000_0001_0000 : 00100
0000_0000_0000_0000_0000_0000_0000_1000 : 00011
0000_0000_0000_0000_0000_0000_0000_0100 : 00010
0000_0000_0000_0000_0000_0000_0000_0010 : 00001
0000_0000_0000_0000_0000_0000_0000_0001 : 00000

Based on this, the minterms are obtained for which the respective output has to be 1.
*/

assign out[4] = |in[31:16];      // continuous assignment statements are used for each individual output bit.

assign out[3] = in[8] | in[9] | in[10] | in[11] | in[12] | in[13] | in[14] | in[15] | 
                in[24] | in[25] | in[26] | in[27] | in[28] | in[29] | in[30] | in[31];

assign out[2] = in[4] | in[5] | in[6] | in[7] | in[12] | in[13] | in[14] | in[15] | 
                in[20] | in[21] | in[22] | in[23] | in[28] | in[29] | in[30] | in[31];

assign out[1] = in[2] | in[3] | in[6] | in[7] | in[10] | in[11] | in[14] | in[15] | 
                in[18] | in[19] | in[22] | in[23] | in[26] | in[27] | in[30] | in[31];

assign out[0] = in[1] | in[3] | in[5] | in[7] | in[9] | in[11] | in[13] | in[15] | 
                in[17] | in[19] | in[21] | in[23] | in[25] | in[27] | in[29] | in[31];
endmodule