// Design a comparator to compare two 16-bit numbers.

module comparator_16(output a_eq_b, a_gr_b, a_ls_b,
                     input [15:0] a, b);

// Easy way to write is as below.
// assign a_eq_b = (a == b);
// assign a_gr_b = (a > b);
// assign a_ls_b = (a < b);
// To consider the work in terms of equations, use the below way

assign a_eq_b = (a[15]~^b[15]) & (a[14]~^b[14]) & (a[13]~^b[13]) & (a[12]~^b[12]) & (a[11]~^b[11]) &
                (a[10]~^b[10]) & (a[9]~^b[9]) & (a[8]~^b[8]) & (a[7]~^b[7]) & (a[6]~^b[6]) &
                (a[5]~^b[5]) & (a[4]~^b[4]) & (a[3]~^b[3]) & (a[2]~^b[2]) & (a[1]~^b[1]) & (a[0]~^b[0]);

assign a_gr_b = (a[15]&(~b[15])) | 
                (a[15]~^b[15])&(a[14]&(~b[14]) |
                (a[14]~^b[14])&(a[13]&(~b[13]) |
                (a[13]~^b[13])&(a[12]&(~b[12]) |
                (a[12]~^b[12])&(a[11]&(~b[11]) |
                (a[11]~^b[11])&(a[10]&(~b[10]) |
                (a[10]~^b[10])&(a[9]&(~b[9]) |
                (a[9]~^b[9])&(a[8]&(~b[8]) |
                (a[8]~^b[8])&(a[7]&(~b[7]) |
                (a[7]~^b[7])&(a[6]&(~b[6]) |
                (a[6]~^b[6])&(a[5]&(~b[5]) |
                (a[5]~^b[5])&(a[4]&(~b[4]) |
                (a[4]~^b[4])&(a[3]&(~b[3]) |
                (a[3]~^b[3])&(a[2]&(~b[2]) |
                (a[2]~^b[2])&(a[1]&(~b[1]) |
                (a[1]~^b[1])&(a[0]&(~b[0])
                )))))))))))))));

assign a_ls_b = (~a[15]&(b[15])) | 
                (a[15]~^b[15])&(~a[14]&(b[14]) |
                (a[14]~^b[14])&(~a[13]&(b[13]) |
                (a[13]~^b[13])&(~a[12]&(b[12]) |
                (a[12]~^b[12])&(~a[11]&(b[11]) |
                (a[11]~^b[11])&(~a[10]&(b[10]) |
                (a[10]~^b[10])&(~a[9]&(b[9]) |
                (a[9]~^b[9])&(~a[8]&(b[8]) |
                (a[8]~^b[8])&(~a[7]&(b[7]) |
                (a[7]~^b[7])&(~a[6]&(b[6]) |
                (a[6]~^b[6])&(~a[5]&(b[5]) |
                (a[5]~^b[5])&(~a[4]&(b[4]) |
                (a[4]~^b[4])&(~a[3]&(b[3]) |
                (a[3]~^b[3])&(~a[2]&(b[2]) |
                (a[2]~^b[2])&(~a[1]&(b[1]) |
                (a[1]~^b[1])&(~a[0]&(b[0])
                )))))))))))))));

endmodule