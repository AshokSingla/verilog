module inverter_not_gate(out, a);
	input a;
	output out;
	assign out = ~a;
endmodule