module buffer(out, a);
	input a;
	output out;
	assign out = a;
endmodule