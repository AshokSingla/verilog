// Design a comparator to compare two 10-bit numbers.

module comparator_10(output a_eq_b, a_ls_b, a_gr_b,
                     input [9:0] a, b);

assign a_eq_b = (a[9]~^b[9]) & (a[8]~^b[8]) & (a[7]~^b[7]) & (a[6]~^b[6]) & (a[5]~^b[5]) &
                (a[4]~^b[4]) & (a[3]~^b[3]) & (a[2]~^b[2]) & (a[1]~^b[1]) & (a[0]~^b[0]) ;

assign a_ls_b = (~a[9] & b[9]) |
                (a[9] & b[9]) & ((~a[8]&b[8]) |
                (a[8] & b[8]) & ((~a[7]&b[7]) |
                (a[7] & b[7]) & ((~a[6]&b[6]) |
                (a[6] & b[6]) & ((~a[5]&b[5]) |
                (a[5] & b[5]) & ((~a[4]&b[4]) |
                (a[4] & b[4]) & ((~a[3]&b[3]) |
                (a[3] & b[3]) & ((~a[2]&b[2]) |
                (a[2] & b[2]) & ((~a[1]&b[1]) |
                (a[1] & b[1]) & ((~a[0]&b[0])
                )))))))));

assign a_gr_b = (a[9] & ~b[9]) |
                (a[9] & b[9]) & ((a[8]&~b[8]) |
                (a[8] & b[8]) & ((a[7]&~b[7]) |
                (a[7] & b[7]) & ((a[6]&~b[6]) |
                (a[6] & b[6]) & ((a[5]&~b[5]) |
                (a[5] & b[5]) & ((a[4]&~b[4]) |
                (a[4] & b[4]) & ((a[3]&~b[3]) |
                (a[3] & b[3]) & ((a[2]&~b[2]) |
                (a[2] & b[2]) & ((a[1]&~b[1]) |
                (a[1] & b[1]) & ((a[0]&~b[0])
                )))))))));                

endmodule                     